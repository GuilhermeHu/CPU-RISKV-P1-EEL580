<?xml version="1.0" encoding="UTF-8" standalone="no"?>
<project source="3.8.0" version="1.0">
  This file is intended to be loaded by Logisim-evolution v3.8.0(https://github.com/logisim-evolution/).

  <lib desc="#Wiring" name="0">
    <tool name="Splitter">
      <a name="facing" val="south"/>
    </tool>
    <tool name="Pin">
      <a name="appearance" val="classic"/>
    </tool>
    <tool name="Probe">
      <a name="appearance" val="classic"/>
      <a name="facing" val="west"/>
    </tool>
    <tool name="Tunnel">
      <a name="facing" val="east"/>
    </tool>
    <tool name="Clock">
      <a name="facing" val="west"/>
    </tool>
    <tool name="Constant">
      <a name="value" val="0x3"/>
      <a name="width" val="2"/>
    </tool>
  </lib>

  <lib desc="#Gates" name="1"/>
  <lib desc="#Plexers" name="2"/>
  <lib desc="#Arithmetic" name="3"/>
  <lib desc="#Memory" name="4"/>
  <lib desc="#I/O" name="5"/>
  <lib desc="#TTL" name="6"/>
  <lib desc="#TCL" name="7"/>
  <lib desc="#Base" name="8"/>
  <lib desc="#BFH-Praktika" name="9"/>
  <lib desc="#Input/Output-Extra" name="10"/>
  <lib desc="#Soc" name="11"/>

  <main name="main"/>
  <options>
    <a name="gateUndefined" val="ignore"/>
    <a name="simlimit" val="1000"/>
    <a name="simrand" val="0"/>
  </options>
  <mappings>
    <tool lib="8" map="Button2" name="Menu Tool"/>
    <tool lib="8" map="Button3" name="Menu Tool"/>
    <tool lib="8" map="Ctrl Button1" name="Menu Tool"/>
  </mappings>
  <toolbar>
    <tool lib="8" name="Poke Tool"/>
    <tool lib="8" name="Edit Tool"/>
    <tool lib="8" name="Wiring Tool"/>
    <tool lib="8" name="Text Tool"/>
    <sep/>
    <tool lib="0" name="Pin"/>
    <tool lib="0" name="Pin">
      <a name="facing" val="west"/>
      <a name="output" val="true"/>
    </tool>
    <sep/>
    <tool lib="1" name="NOT Gate"/>
    <tool lib="1" name="AND Gate"/>
    <tool lib="1" name="OR Gate"/>
    <tool lib="1" name="XOR Gate"/>
    <tool lib="1" name="NAND Gate"/>
    <tool lib="1" name="NOR Gate"/>
    <sep/>
    <tool lib="4" name="D Flip-Flop"/>
    <tool lib="4" name="Register"/>
  </toolbar>
  <circuit name="main">
    <a name="appearance" val="logisim_evolution"/>
    <a name="circuit" val="main"/>
    <a name="circuitnamedboxfixedsize" val="true"/>
    <a name="simulationFrequency" val="1.0"/>
    <comp lib="0" loc="(1020,560)" name="Splitter">
      <a name="appear" val="right"/>
      <a name="fanout" val="32"/>
      <a name="incoming" val="32"/>
    </comp>
    <comp lib="0" loc="(1110,1060)" name="Probe">
      <a name="appearance" val="classic"/>
    </comp>
    <comp lib="0" loc="(1110,690)" name="Splitter">
      <a name="appear" val="right"/>
      <a name="facing" val="west"/>
      <a name="fanout" val="5"/>
      <a name="incoming" val="5"/>
    </comp>
    <comp lib="0" loc="(1110,710)" name="Splitter">
      <a name="facing" val="west"/>
      <a name="fanout" val="5"/>
      <a name="incoming" val="5"/>
    </comp>
    <comp lib="0" loc="(1110,830)" name="Splitter">
      <a name="facing" val="west"/>
      <a name="fanout" val="4"/>
      <a name="incoming" val="4"/>
    </comp>
    <comp lib="0" loc="(1120,760)" name="Splitter">
      <a name="facing" val="west"/>
      <a name="fanout" val="5"/>
      <a name="incoming" val="5"/>
    </comp>
    <comp lib="0" loc="(1130,640)" name="Splitter">
      <a name="appear" val="right"/>
      <a name="facing" val="west"/>
      <a name="fanout" val="7"/>
      <a name="incoming" val="7"/>
    </comp>
    <comp lib="0" loc="(1150,450)" name="Pin">
      <a name="appearance" val="NewPins"/>
      <a name="width" val="5"/>
    </comp>
    <comp lib="0" loc="(120,420)" name="Constant">
      <a name="value" val="0x0"/>
    </comp>
    <comp lib="0" loc="(130,610)" name="Pin">
      <a name="appearance" val="NewPins"/>
      <a name="facing" val="south"/>
    </comp>
    <comp lib="0" loc="(1390,440)" name="Probe">
      <a name="appearance" val="classic"/>
    </comp>
    <comp lib="0" loc="(1510,1190)" name="Splitter">
      <a name="appear" val="right"/>
    </comp>
    <comp lib="0" loc="(1520,1170)" name="Splitter">
      <a name="appear" val="right"/>
    </comp>
    <comp lib="0" loc="(1570,1040)" name="Splitter">
      <a name="facing" val="west"/>
      <a name="fanout" val="6"/>
      <a name="incoming" val="6"/>
      <a name="spacing" val="2"/>
    </comp>
    <comp lib="0" loc="(1630,980)" name="Splitter">
      <a name="facing" val="west"/>
      <a name="fanout" val="4"/>
      <a name="incoming" val="4"/>
      <a name="spacing" val="2"/>
    </comp>
    <comp lib="0" loc="(1650,1090)" name="Splitter">
      <a name="facing" val="west"/>
      <a name="fanout" val="3"/>
      <a name="incoming" val="3"/>
      <a name="spacing" val="2"/>
    </comp>
    <comp lib="0" loc="(1700,1080)" name="Constant">
      <a name="value" val="0x0"/>
      <a name="width" val="3"/>
    </comp>
    <comp lib="0" loc="(1700,920)" name="Constant">
      <a name="value" val="0x0"/>
      <a name="width" val="6"/>
    </comp>
    <comp lib="0" loc="(1700,990)" name="Constant">
      <a name="value" val="0x0"/>
      <a name="width" val="4"/>
    </comp>
    <comp lib="0" loc="(1900,200)" name="Splitter">
      <a name="appear" val="right"/>
    </comp>
    <comp lib="0" loc="(1910,680)" name="Splitter">
      <a name="appear" val="right"/>
      <a name="fanout" val="4"/>
      <a name="incoming" val="4"/>
    </comp>
    <comp lib="0" loc="(1920,1150)" name="Splitter">
      <a name="facing" val="west"/>
      <a name="fanout" val="6"/>
      <a name="incoming" val="6"/>
      <a name="spacing" val="2"/>
    </comp>
    <comp lib="0" loc="(1950,730)" name="Splitter">
      <a name="appear" val="right"/>
      <a name="facing" val="west"/>
    </comp>
    <comp lib="0" loc="(2030,440)" name="Constant">
      <a name="value" val="0x0"/>
      <a name="width" val="32"/>
    </comp>
    <comp lib="0" loc="(250,840)" name="Splitter">
      <a name="appear" val="right"/>
      <a name="fanout" val="8"/>
      <a name="incoming" val="8"/>
    </comp>
    <comp lib="0" loc="(2760,610)" name="Splitter">
      <a name="appear" val="right"/>
      <a name="fanout" val="6"/>
      <a name="incoming" val="6"/>
      <a name="spacing" val="2"/>
    </comp>
    <comp lib="0" loc="(2850,1020)" name="Splitter">
      <a name="facing" val="west"/>
      <a name="fanout" val="3"/>
      <a name="incoming" val="3"/>
    </comp>
    <comp lib="0" loc="(2960,640)" name="Splitter">
      <a name="appear" val="right"/>
      <a name="fanout" val="32"/>
      <a name="incoming" val="32"/>
    </comp>
    <comp lib="0" loc="(3010,640)" name="Splitter">
      <a name="facing" val="west"/>
      <a name="fanout" val="24"/>
      <a name="incoming" val="24"/>
    </comp>
    <comp lib="0" loc="(3620,570)" name="Splitter">
      <a name="appear" val="right"/>
      <a name="fanout" val="3"/>
      <a name="incoming" val="3"/>
    </comp>
    <comp lib="0" loc="(3710,570)" name="Splitter">
      <a name="facing" val="west"/>
    </comp>
    <comp lib="0" loc="(430,600)" name="Splitter">
      <a name="appear" val="right"/>
      <a name="fanout" val="32"/>
      <a name="incoming" val="32"/>
    </comp>
    <comp lib="0" loc="(470,600)" name="Splitter">
      <a name="facing" val="west"/>
      <a name="fanout" val="24"/>
      <a name="incoming" val="24"/>
    </comp>
    <comp lib="0" loc="(500,310)" name="Constant">
      <a name="width" val="32"/>
    </comp>
    <comp lib="0" loc="(70,870)" name="Clock"/>
    <comp lib="1" loc="(2900,400)" name="OR Gate">
      <a name="size" val="30"/>
    </comp>
    <comp lib="1" loc="(2910,270)" name="OR Gate">
      <a name="facing" val="north"/>
    </comp>
    <comp lib="1" loc="(2930,330)" name="AND Gate">
      <a name="facing" val="north"/>
    </comp>
    <comp lib="1" loc="(2960,460)" name="NOT Gate">
      <a name="facing" val="north"/>
    </comp>
    <comp lib="2" loc="(1550,180)" name="Multiplexer">
      <a name="facing" val="north"/>
      <a name="select" val="2"/>
      <a name="selloc" val="tr"/>
      <a name="width" val="32"/>
    </comp>
    <comp lib="2" loc="(1760,1070)" name="Multiplexer">
      <a name="width" val="3"/>
    </comp>
    <comp lib="2" loc="(1760,910)" name="Multiplexer">
      <a name="width" val="6"/>
    </comp>
    <comp lib="2" loc="(1760,980)" name="Multiplexer">
      <a name="width" val="4"/>
    </comp>
    <comp lib="2" loc="(2080,560)" name="Multiplexer">
      <a name="width" val="32"/>
    </comp>
    <comp lib="2" loc="(2100,620)" name="Multiplexer">
      <a name="width" val="32"/>
    </comp>
    <comp lib="2" loc="(2120,790)" name="Multiplexer">
      <a name="select" val="2"/>
      <a name="width" val="32"/>
    </comp>
    <comp lib="2" loc="(2180,750)" name="Multiplexer">
      <a name="select" val="2"/>
      <a name="width" val="32"/>
    </comp>
    <comp lib="2" loc="(2950,420)" name="Multiplexer">
      <a name="facing" val="north"/>
    </comp>
    <comp lib="2" loc="(3730,540)" name="Multiplexer">
      <a name="select" val="2"/>
      <a name="width" val="32"/>
    </comp>
    <comp lib="2" loc="(80,400)" name="Multiplexer">
      <a name="facing" val="south"/>
      <a name="selloc" val="tr"/>
      <a name="width" val="32"/>
    </comp>
    <comp lib="4" loc="(130,410)" name="D Flip-Flop">
      <a name="appearance" val="logisim_evolution"/>
    </comp>
    <comp lib="4" loc="(250,840)" name="Counter">
      <a name="appearance" val="classic"/>
    </comp>
    <comp lib="4" loc="(3090,630)" name="RAM">
      <a name="addrWidth" val="24"/>
      <a name="appearance" val="logisim_evolution"/>
      <a name="dataWidth" val="32"/>
    </comp>
    <comp lib="4" loc="(480,590)" name="ROM">
      <a name="addrWidth" val="24"/>
      <a name="appearance" val="logisim_evolution"/>
      <a name="contents">addr/data: 24 32                     -- Respectivamente, largura do enedereço e e largura dos dados, em bits
9563  -- Valor que é armazenado no endereço inicial da ROM
</a>                                                            -- SEGUNDO O CHAT GPT, PODEMOS MUDAR ESSAS DUAS LINHAS PRA CIMA
      <a name="dataWidth" val="32"/>
      <a name="labelvisible" val="true"/>
    </comp>
    <comp loc="(1160,1320)" name="Harzard">
      <a name="appearance" val="logisim_evolution"/>
    </comp>
    <comp loc="(1470,560)" name="register_file">
      <a name="appearance" val="logisim_evolution"/>
    </comp>
    <comp loc="(1470,910)" name="ImmGen">
      <a name="appearance" val="logisim_evolution"/>
    </comp>
    <comp loc="(1470,990)" name="Control_Unit">
      <a name="appearance" val="logisim_evolution"/>
    </comp>
    <comp loc="(1880,520)" name="IDEX">
      <a name="appearance" val="logisim_evolution"/>
    </comp>
    <comp loc="(2380,510)" name="somador">
      <a name="appearance" val="logisim_evolution"/>
    </comp>
    <comp loc="(2430,600)" name="ALU">
      <a name="appearance" val="logisim_evolution"/>
    </comp>
    <comp loc="(2430,850)" name="ALU_Control">
      <a name="appearance" val="logisim_evolution"/>
    </comp>
    <comp loc="(2570,1130)" name="Forward">
      <a name="appearance" val="logisim_evolution"/>
    </comp>
    <comp loc="(2750,490)" name="EXMEM">
      <a name="appearance" val="logisim_evolution"/>
    </comp>
    <comp loc="(3600,510)" name="MEMWB">
      <a name="appearance" val="logisim_evolution"/>
    </comp>
    <comp loc="(420,600)" name="PC2">
      <a name="appearance" val="logisim_evolution"/>
    </comp>
    <comp loc="(720,290)" name="somador">
      <a name="appearance" val="logisim_evolution"/>
      <a name="labelvisible" val="true"/>
    </comp>
    <comp loc="(980,540)" name="IFID">
      <a name="appearance" val="logisim_evolution"/>
    </comp>

    <wire from="(100,380)" to="(210,380)"/>
    <wire from="(100,460)" to="(100,870)"/>
    <wire from="(100,460)" to="(120,460)"/>
    <wire from="(100,870)" to="(190,870)"/>
    <wire from="(1000,580)" to="(1000,910)"/>
    <wire from="(1000,580)" to="(1020,580)"/>
    <wire from="(1000,910)" to="(1070,910)"/>
    <wire from="(1020,560)" to="(1020,580)"/>
    <wire from="(1040,570)" to="(1110,570)"/>
    <wire from="(1040,580)" to="(1110,580)"/>
    <wire from="(1040,590)" to="(1110,590)"/>
    <wire from="(1040,600)" to="(1110,600)"/>
    <wire from="(1040,610)" to="(1110,610)"/>
    <wire from="(1040,620)" to="(1110,620)"/>
    <wire from="(1040,630)" to="(1110,630)"/>
    <wire from="(1040,640)" to="(1090,640)"/>
    <wire from="(1040,650)" to="(1090,650)"/>
    <wire from="(1040,660)" to="(1090,660)"/>
    <wire from="(1040,670)" to="(1090,670)"/>
    <wire from="(1040,680)" to="(1090,680)"/>
    <wire from="(1040,690)" to="(1070,690)"/>
    <wire from="(1040,700)" to="(1060,700)"/>
    <wire from="(1040,710)" to="(1050,710)"/>
    <wire from="(1040,720)" to="(1090,720)"/>
    <wire from="(1040,730)" to="(1090,730)"/>
    <wire from="(1040,740)" to="(1090,740)"/>
    <wire from="(1040,750)" to="(1090,750)"/>
    <wire from="(1040,760)" to="(1090,760)"/>
    <wire from="(1040,770)" to="(1100,770)"/>
    <wire from="(1040,780)" to="(1100,780)"/>
    <wire from="(1040,790)" to="(1100,790)"/>
    <wire from="(1040,800)" to="(1100,800)"/>
    <wire from="(1040,810)" to="(1100,810)"/>
    <wire from="(1040,870)" to="(1090,870)"/>
    <wire from="(1050,710)" to="(1050,860)"/>
    <wire from="(1050,860)" to="(1090,860)"/>
    <wire from="(1060,700)" to="(1060,850)"/>
    <wire from="(1060,850)" to="(1090,850)"/>
    <wire from="(1070,1010)" to="(1120,1010)"/>
    <wire from="(1070,690)" to="(1070,840)"/>
    <wire from="(1070,840)" to="(1090,840)"/>
    <wire from="(1070,910)" to="(1070,1010)"/>
    <wire from="(1070,910)" to="(1250,910)"/>
    <wire from="(1110,1060)" to="(1120,1060)"/>
    <wire from="(1110,690)" to="(1180,690)"/>
    <wire from="(1110,710)" to="(1160,710)"/>
    <wire from="(1110,830)" to="(1580,830)"/>
    <wire from="(1120,1010)" to="(1120,1060)"/>
    <wire from="(1120,760)" to="(1170,760)"/>
    <wire from="(1130,640)" to="(1130,990)"/>
    <wire from="(1130,990)" to="(1250,990)"/>
    <wire from="(1150,450)" to="(1170,450)"/>
    <wire from="(1160,1320)" to="(1170,1320)"/>
    <wire from="(1160,620)" to="(1160,710)"/>
    <wire from="(1160,620)" to="(1250,620)"/>
    <wire from="(1160,710)" to="(1160,740)"/>
    <wire from="(1160,740)" to="(1160,1150)"/>
    <wire from="(1160,740)" to="(1660,740)"/>
    <wire from="(1170,1300)" to="(1170,1320)"/>
    <wire from="(1170,1300)" to="(1710,1300)"/>
    <wire from="(1170,450)" to="(1170,580)"/>
    <wire from="(1170,580)" to="(1250,580)"/>
    <wire from="(1170,640)" to="(1170,760)"/>
    <wire from="(1170,640)" to="(1250,640)"/>
    <wire from="(1170,760)" to="(1170,1160)"/>
    <wire from="(1170,760)" to="(1660,760)"/>
    <wire from="(1180,690)" to="(1180,730)"/>
    <wire from="(1180,730)" to="(1500,730)"/>
    <wire from="(1190,1410)" to="(2130,1410)"/>
    <wire from="(1190,560)" to="(1190,1410)"/>
    <wire from="(1190,560)" to="(1250,560)"/>
    <wire from="(1210,1400)" to="(3690,1400)"/>
    <wire from="(1210,600)" to="(1210,1400)"/>
    <wire from="(1210,600)" to="(1250,600)"/>
    <wire from="(1220,1380)" to="(2300,1380)"/>
    <wire from="(1220,660)" to="(1220,1380)"/>
    <wire from="(1220,660)" to="(1250,660)"/>
    <wire from="(1240,1460)" to="(2240,1460)"/>
    <wire from="(1240,680)" to="(1240,1460)"/>
    <wire from="(1240,680)" to="(1250,680)"/>
    <wire from="(130,1300)" to="(750,1300)"/>
    <wire from="(130,610)" to="(130,620)"/>
    <wire from="(130,620)" to="(200,620)"/>
    <wire from="(130,660)" to="(130,1300)"/>
    <wire from="(130,660)" to="(200,660)"/>
    <wire from="(1390,440)" to="(1480,440)"/>
    <wire from="(1470,1010)" to="(1610,1010)"/>
    <wire from="(1470,1030)" to="(1500,1030)"/>
    <wire from="(1470,1050)" to="(1550,1050)"/>
    <wire from="(1470,1070)" to="(1550,1070)"/>
    <wire from="(1470,1090)" to="(1550,1090)"/>
    <wire from="(1470,1110)" to="(1550,1110)"/>
    <wire from="(1470,1130)" to="(1550,1130)"/>
    <wire from="(1470,1150)" to="(1550,1150)"/>
    <wire from="(1470,1170)" to="(1520,1170)"/>
    <wire from="(1470,1190)" to="(1510,1190)"/>
    <wire from="(1470,560)" to="(1660,560)"/>
    <wire from="(1470,580)" to="(1660,580)"/>
    <wire from="(1470,600)" to="(1480,600)"/>
    <wire from="(1470,910)" to="(1540,910)"/>
    <wire from="(1470,990)" to="(1610,990)"/>
    <wire from="(1480,440)" to="(1480,600)"/>
    <wire from="(150,600)" to="(150,780)"/>
    <wire from="(150,600)" to="(190,600)"/>
    <wire from="(150,780)" to="(300,780)"/>
    <wire from="(1500,1030)" to="(1500,1220)"/>
    <wire from="(1500,1220)" to="(1630,1220)"/>
    <wire from="(1500,640)" to="(1500,730)"/>
    <wire from="(1500,640)" to="(1660,640)"/>
    <wire from="(1530,1200)" to="(1610,1200)"/>
    <wire from="(1530,1210)" to="(1620,1210)"/>
    <wire from="(1530,220)" to="(1530,290)"/>
    <wire from="(1540,1180)" to="(1590,1180)"/>
    <wire from="(1540,1190)" to="(1600,1190)"/>
    <wire from="(1540,220)" to="(1540,290)"/>
    <wire from="(1540,290)" to="(2800,290)"/>
    <wire from="(1540,600)" to="(1540,910)"/>
    <wire from="(1540,600)" to="(1660,600)"/>
    <wire from="(1550,150)" to="(1550,180)"/>
    <wire from="(1550,220)" to="(1550,270)"/>
    <wire from="(1550,270)" to="(1790,270)"/>
    <wire from="(1560,220)" to="(1560,250)"/>
    <wire from="(1560,250)" to="(1790,250)"/>
    <wire from="(1570,200)" to="(1900,200)"/>
    <wire from="(1570,900)" to="(1570,1040)"/>
    <wire from="(1570,900)" to="(1730,900)"/>
    <wire from="(1580,620)" to="(1580,830)"/>
    <wire from="(1580,620)" to="(1660,620)"/>
    <wire from="(1590,1030)" to="(1590,1180)"/>
    <wire from="(1590,1030)" to="(1610,1030)"/>
    <wire from="(1590,660)" to="(1590,850)"/>
    <wire from="(1590,660)" to="(1660,660)"/>
    <wire from="(1590,850)" to="(1820,850)"/>
    <wire from="(1600,1050)" to="(1600,1190)"/>
    <wire from="(1600,1050)" to="(1610,1050)"/>
    <wire from="(1600,680)" to="(1600,870)"/>
    <wire from="(1600,680)" to="(1660,680)"/>
    <wire from="(1600,870)" to="(1790,870)"/>
    <wire from="(1610,1100)" to="(1610,1200)"/>
    <wire from="(1610,1100)" to="(1630,1100)"/>
    <wire from="(1610,700)" to="(1610,860)"/>
    <wire from="(1610,700)" to="(1660,700)"/>
    <wire from="(1610,860)" to="(1810,860)"/>
    <wire from="(1620,1120)" to="(1620,1210)"/>
    <wire from="(1620,1120)" to="(1630,1120)"/>
    <wire from="(1620,720)" to="(1620,890)"/>
    <wire from="(1620,720)" to="(1660,720)"/>
    <wire from="(1630,1140)" to="(1630,1220)"/>
    <wire from="(1630,970)" to="(1630,980)"/>
    <wire from="(1630,970)" to="(1730,970)"/>
    <wire from="(1640,490)" to="(1640,520)"/>
    <wire from="(1640,490)" to="(2520,490)"/>
    <wire from="(1640,520)" to="(1660,520)"/>
    <wire from="(1650,1060)" to="(1650,1090)"/>
    <wire from="(1650,1060)" to="(1730,1060)"/>
    <wire from="(1700,1080)" to="(1730,1080)"/>
    <wire from="(1700,920)" to="(1730,920)"/>
    <wire from="(1700,990)" to="(1730,990)"/>
    <wire from="(1710,1010)" to="(1710,1100)"/>
    <wire from="(1710,1010)" to="(1740,1010)"/>
    <wire from="(1710,1100)" to="(1710,1300)"/>
    <wire from="(1710,1100)" to="(1740,1100)"/>
    <wire from="(1710,940)" to="(1710,1010)"/>
    <wire from="(1710,940)" to="(1740,940)"/>
    <wire from="(1740,1000)" to="(1740,1010)"/>
    <wire from="(1740,1090)" to="(1740,1100)"/>
    <wire from="(1740,930)" to="(1740,940)"/>
    <wire from="(1760,1070)" to="(1820,1070)"/>
    <wire from="(1760,910)" to="(1790,910)"/>
    <wire from="(1760,980)" to="(1810,980)"/>
    <wire from="(1790,140)" to="(1790,250)"/>
    <wire from="(1790,140)" to="(3030,140)"/>
    <wire from="(1790,250)" to="(1790,270)"/>
    <wire from="(1790,870)" to="(1790,910)"/>
    <wire from="(180,420)" to="(210,420)"/>
    <wire from="(1810,860)" to="(1810,980)"/>
    <wire from="(1820,850)" to="(1820,1070)"/>
    <wire from="(1880,1100)" to="(2200,1100)"/>
    <wire from="(1880,520)" to="(2010,520)"/>
    <wire from="(1880,540)" to="(1950,540)"/>
    <wire from="(1880,560)" to="(2000,560)"/>
    <wire from="(1880,580)" to="(2030,580)"/>
    <wire from="(1880,600)" to="(2020,600)"/>
    <wire from="(1880,620)" to="(1990,620)"/>
    <wire from="(1880,640)" to="(1980,640)"/>
    <wire from="(1880,660)" to="(1970,660)"/>
    <wire from="(1880,680)" to="(1910,680)"/>
    <wire from="(1880,700)" to="(1910,700)"/>
    <wire from="(1880,720)" to="(1900,720)"/>
    <wire from="(1880,740)" to="(1880,1100)"/>
    <wire from="(1890,1160)" to="(1890,1250)"/>
    <wire from="(1890,1160)" to="(1900,1160)"/>
    <wire from="(190,1460)" to="(830,1460)"/>
    <wire from="(190,540)" to="(190,600)"/>
    <wire from="(190,540)" to="(750,540)"/>
    <wire from="(190,600)" to="(200,600)"/>
    <wire from="(190,870)" to="(190,1460)"/>
    <wire from="(190,870)" to="(230,870)"/>
    <wire from="(1900,1080)" to="(2220,1080)"/>
    <wire from="(1900,720)" to="(1900,1080)"/>
    <wire from="(1910,700)" to="(1910,950)"/>
    <wire from="(1910,950)" to="(2510,950)"/>
    <wire from="(1920,1150)" to="(1970,1150)"/>
    <wire from="(1920,210)" to="(2910,210)"/>
    <wire from="(1920,220)" to="(2840,220)"/>
    <wire from="(1930,690)" to="(2080,690)"/>
    <wire from="(1930,700)" to="(2060,700)"/>
    <wire from="(1950,540)" to="(1950,550)"/>
    <wire from="(1950,550)" to="(2050,550)"/>
    <wire from="(1950,730)" to="(1960,730)"/>
    <wire from="(1960,730)" to="(1960,870)"/>
    <wire from="(1960,870)" to="(2210,870)"/>
    <wire from="(1970,660)" to="(1970,940)"/>
    <wire from="(1970,940)" to="(1970,1150)"/>
    <wire from="(1970,940)" to="(2490,940)"/>
    <wire from="(1980,640)" to="(1980,930)"/>
    <wire from="(1980,930)" to="(2480,930)"/>
    <wire from="(1990,620)" to="(1990,920)"/>
    <wire from="(1990,920)" to="(1990,1280)"/>
    <wire from="(1990,920)" to="(2470,920)"/>
    <wire from="(2000,560)" to="(2000,610)"/>
    <wire from="(2000,610)" to="(2000,910)"/>
    <wire from="(2000,610)" to="(2070,610)"/>
    <wire from="(2000,910)" to="(2460,910)"/>
    <wire from="(2010,510)" to="(2010,520)"/>
    <wire from="(2010,510)" to="(2160,510)"/>
    <wire from="(2020,600)" to="(2020,850)"/>
    <wire from="(2020,850)" to="(2210,850)"/>
    <wire from="(2030,440)" to="(2040,440)"/>
    <wire from="(2030,530)" to="(2030,580)"/>
    <wire from="(2030,530)" to="(2160,530)"/>
    <wire from="(2030,580)" to="(2030,630)"/>
    <wire from="(2030,630)" to="(2070,630)"/>
    <wire from="(2040,440)" to="(2040,570)"/>
    <wire from="(2040,570)" to="(2050,570)"/>
    <wire from="(2050,1060)" to="(2920,1060)"/>
    <wire from="(2050,750)" to="(2050,790)"/>
    <wire from="(2050,750)" to="(2140,750)"/>
    <wire from="(2050,790)" to="(2050,1060)"/>
    <wire from="(2050,790)" to="(2080,790)"/>
    <wire from="(2060,1040)" to="(2130,1040)"/>
    <wire from="(2060,580)" to="(2060,700)"/>
    <wire from="(2060,780)" to="(2060,1040)"/>
    <wire from="(2060,780)" to="(2080,780)"/>
    <wire from="(2070,740)" to="(2070,770)"/>
    <wire from="(2070,740)" to="(2110,740)"/>
    <wire from="(2070,770)" to="(2080,770)"/>
    <wire from="(2080,560)" to="(2120,560)"/>
    <wire from="(2080,640)" to="(2080,690)"/>
    <wire from="(210,380)" to="(210,420)"/>
    <wire from="(2100,620)" to="(2110,620)"/>
    <wire from="(2100,810)" to="(2100,990)"/>
    <wire from="(2100,990)" to="(2600,990)"/>
    <wire from="(2110,620)" to="(2110,740)"/>
    <wire from="(2120,560)" to="(2120,730)"/>
    <wire from="(2120,730)" to="(2140,730)"/>
    <wire from="(2120,790)" to="(2210,790)"/>
    <wire from="(2130,1040)" to="(2130,1410)"/>
    <wire from="(2130,1410)" to="(3740,1410)"/>
    <wire from="(2130,740)" to="(2130,1040)"/>
    <wire from="(2130,740)" to="(2140,740)"/>
    <wire from="(2160,600)" to="(2160,720)"/>
    <wire from="(2160,600)" to="(2210,600)"/>
    <wire from="(2160,720)" to="(2190,720)"/>
    <wire from="(2160,770)" to="(2160,970)"/>
    <wire from="(2160,970)" to="(2570,970)"/>
    <wire from="(2180,620)" to="(2180,700)"/>
    <wire from="(2180,620)" to="(2210,620)"/>
    <wire from="(2180,700)" to="(2210,700)"/>
    <wire from="(2180,750)" to="(2190,750)"/>
    <wire from="(2190,720)" to="(2190,750)"/>
    <wire from="(2200,1100)" to="(2200,1210)"/>
    <wire from="(2200,1210)" to="(2350,1210)"/>
    <wire from="(2200,640)" to="(2200,680)"/>
    <wire from="(2200,640)" to="(2210,640)"/>
    <wire from="(2200,680)" to="(2440,680)"/>
    <wire from="(2210,700)" to="(2210,790)"/>
    <wire from="(2220,1080)" to="(2220,1190)"/>
    <wire from="(2220,1190)" to="(2350,1190)"/>
    <wire from="(2240,1130)" to="(2240,1460)"/>
    <wire from="(2240,1130)" to="(2350,1130)"/>
    <wire from="(2240,1460)" to="(3050,1460)"/>
    <wire from="(230,860)" to="(230,870)"/>
    <wire from="(2300,1230)" to="(2300,1380)"/>
    <wire from="(2300,1230)" to="(2350,1230)"/>
    <wire from="(2300,1380)" to="(3650,1380)"/>
    <wire from="(2320,1030)" to="(2320,1170)"/>
    <wire from="(2320,1030)" to="(2830,1030)"/>
    <wire from="(2320,1170)" to="(2350,1170)"/>
    <wire from="(2330,1100)" to="(2330,1150)"/>
    <wire from="(2330,1100)" to="(3680,1100)"/>
    <wire from="(2330,1150)" to="(2350,1150)"/>
    <wire from="(2330,1250)" to="(2330,1290)"/>
    <wire from="(2330,1250)" to="(2350,1250)"/>
    <wire from="(2330,1290)" to="(3030,1290)"/>
    <wire from="(2380,510)" to="(2530,510)"/>
    <wire from="(240,860)" to="(240,890)"/>
    <wire from="(2430,600)" to="(2440,600)"/>
    <wire from="(2430,620)" to="(2450,620)"/>
    <wire from="(2430,850)" to="(2440,850)"/>
    <wire from="(2440,550)" to="(2440,600)"/>
    <wire from="(2440,550)" to="(2530,550)"/>
    <wire from="(2440,680)" to="(2440,850)"/>
    <wire from="(2450,530)" to="(2450,620)"/>
    <wire from="(2450,530)" to="(2530,530)"/>
    <wire from="(2460,570)" to="(2460,910)"/>
    <wire from="(2460,570)" to="(2530,570)"/>
    <wire from="(2470,590)" to="(2470,920)"/>
    <wire from="(2470,590)" to="(2530,590)"/>
    <wire from="(2480,610)" to="(2480,930)"/>
    <wire from="(2480,610)" to="(2530,610)"/>
    <wire from="(2490,630)" to="(2490,940)"/>
    <wire from="(2490,630)" to="(2530,630)"/>
    <wire from="(2510,650)" to="(2510,950)"/>
    <wire from="(2510,650)" to="(2530,650)"/>
    <wire from="(2520,240)" to="(2520,490)"/>
    <wire from="(2520,240)" to="(3340,240)"/>
    <wire from="(2520,490)" to="(2530,490)"/>
    <wire from="(2570,1150)" to="(2600,1150)"/>
    <wire from="(2570,970)" to="(2570,1130)"/>
    <wire from="(2600,990)" to="(2600,1150)"/>
    <wire from="(270,850)" to="(300,850)"/>
    <wire from="(2750,1370)" to="(3360,1370)"/>
    <wire from="(2750,490)" to="(2800,490)"/>
    <wire from="(2750,510)" to="(2940,510)"/>
    <wire from="(2750,530)" to="(2920,530)"/>
    <wire from="(2750,550)" to="(2890,550)"/>
    <wire from="(2750,570)" to="(3030,570)"/>
    <wire from="(2750,590)" to="(2910,590)"/>
    <wire from="(2750,610)" to="(2760,610)"/>
    <wire from="(2750,630)" to="(2750,1370)"/>
    <wire from="(2780,620)" to="(2880,620)"/>
    <wire from="(2780,640)" to="(2870,640)"/>
    <wire from="(2780,660)" to="(2790,660)"/>
    <wire from="(2780,680)" to="(2830,680)"/>
    <wire from="(2780,700)" to="(2810,700)"/>
    <wire from="(2780,720)" to="(2840,720)"/>
    <wire from="(2790,390)" to="(2790,660)"/>
    <wire from="(2790,390)" to="(2870,390)"/>
    <wire from="(2800,250)" to="(2800,290)"/>
    <wire from="(2800,250)" to="(3270,250)"/>
    <wire from="(2800,290)" to="(2800,490)"/>
    <wire from="(2810,330)" to="(2810,700)"/>
    <wire from="(2810,330)" to="(2890,330)"/>
    <wire from="(2830,440)" to="(2830,680)"/>
    <wire from="(2830,440)" to="(2850,440)"/>
    <wire from="(2840,220)" to="(2840,720)"/>
    <wire from="(2850,1020)" to="(2910,1020)"/>
    <wire from="(2850,410)" to="(2850,440)"/>
    <wire from="(2850,410)" to="(2870,410)"/>
    <wire from="(2850,440)" to="(2930,440)"/>
    <wire from="(2870,640)" to="(2870,990)"/>
    <wire from="(2870,990)" to="(3010,990)"/>
    <wire from="(2880,620)" to="(2880,980)"/>
    <wire from="(2880,980)" to="(3020,980)"/>
    <wire from="(2890,320)" to="(2890,330)"/>
    <wire from="(2890,550)" to="(2890,970)"/>
    <wire from="(2890,970)" to="(3090,970)"/>
    <wire from="(2900,400)" to="(2910,400)"/>
    <wire from="(2910,210)" to="(2910,270)"/>
    <wire from="(2910,380)" to="(2910,400)"/>
    <wire from="(2910,590)" to="(2910,1020)"/>
    <wire from="(2910,590)" to="(3380,590)"/>
    <wire from="(2920,530)" to="(2920,640)"/>
    <wire from="(2920,530)" to="(3030,530)"/>
    <wire from="(2920,640)" to="(2920,1060)"/>
    <wire from="(2920,640)" to="(2960,640)"/>
    <wire from="(2930,320)" to="(2930,330)"/>
    <wire from="(2940,450)" to="(2940,510)"/>
    <wire from="(2940,510)" to="(2960,510)"/>
    <wire from="(2950,380)" to="(2950,420)"/>
    <wire from="(2960,450)" to="(2960,460)"/>
    <wire from="(2960,490)" to="(2960,510)"/>
    <wire from="(2980,650)" to="(2990,650)"/>
    <wire from="(2980,660)" to="(2990,660)"/>
    <wire from="(2980,670)" to="(2990,670)"/>
    <wire from="(2980,680)" to="(2990,680)"/>
    <wire from="(2980,690)" to="(2990,690)"/>
    <wire from="(2980,700)" to="(2990,700)"/>
    <wire from="(2980,710)" to="(2990,710)"/>
    <wire from="(2980,720)" to="(2990,720)"/>
    <wire from="(2980,730)" to="(2990,730)"/>
    <wire from="(2980,740)" to="(2990,740)"/>
    <wire from="(2980,750)" to="(2990,750)"/>
    <wire from="(2980,760)" to="(2990,760)"/>
    <wire from="(2980,770)" to="(2990,770)"/>
    <wire from="(2980,780)" to="(2990,780)"/>
    <wire from="(2980,790)" to="(2990,790)"/>
    <wire from="(2980,800)" to="(2990,800)"/>
    <wire from="(2980,810)" to="(2990,810)"/>
    <wire from="(2980,820)" to="(2990,820)"/>
    <wire from="(2980,830)" to="(2990,830)"/>
    <wire from="(2980,840)" to="(2990,840)"/>
    <wire from="(2980,850)" to="(2990,850)"/>
    <wire from="(2980,860)" to="(2990,860)"/>
    <wire from="(2980,870)" to="(2990,870)"/>
    <wire from="(2980,880)" to="(2990,880)"/>
    <wire from="(300,780)" to="(300,850)"/>
    <wire from="(3010,640)" to="(3090,640)"/>
    <wire from="(3010,680)" to="(3010,990)"/>
    <wire from="(3010,680)" to="(3090,680)"/>
    <wire from="(3020,690)" to="(3020,980)"/>
    <wire from="(3020,690)" to="(3090,690)"/>
    <wire from="(3030,140)" to="(3030,530)"/>
    <wire from="(3030,530)" to="(3030,550)"/>
    <wire from="(3030,550)" to="(3380,550)"/>
    <wire from="(3030,570)" to="(3030,1290)"/>
    <wire from="(3030,570)" to="(3380,570)"/>
    <wire from="(3050,700)" to="(3050,1460)"/>
    <wire from="(3050,700)" to="(3090,700)"/>
    <wire from="(3090,720)" to="(3090,970)"/>
    <wire from="(3270,250)" to="(3270,620)"/>
    <wire from="(3270,620)" to="(3380,620)"/>
    <wire from="(3330,720)" to="(3340,720)"/>
    <wire from="(3340,240)" to="(3340,510)"/>
    <wire from="(3340,510)" to="(3380,510)"/>
    <wire from="(3340,530)" to="(3340,720)"/>
    <wire from="(3340,530)" to="(3380,530)"/>
    <wire from="(3360,610)" to="(3360,1370)"/>
    <wire from="(3360,610)" to="(3380,610)"/>
    <wire from="(3380,620)" to="(3380,630)"/>
    <wire from="(3600,510)" to="(3650,510)"/>
    <wire from="(3600,530)" to="(3630,530)"/>
    <wire from="(3600,550)" to="(3650,550)"/>
    <wire from="(3600,570)" to="(3620,570)"/>
    <wire from="(3600,590)" to="(3610,590)"/>
    <wire from="(3600,610)" to="(3600,640)"/>
    <wire from="(3600,640)" to="(3670,640)"/>
    <wire from="(3610,590)" to="(3610,610)"/>
    <wire from="(3610,610)" to="(3660,610)"/>
    <wire from="(3630,520)" to="(3630,530)"/>
    <wire from="(3630,520)" to="(3690,520)"/>
    <wire from="(3640,580)" to="(3680,580)"/>
    <wire from="(3640,590)" to="(3690,590)"/>
    <wire from="(3640,600)" to="(3690,600)"/>
    <wire from="(3650,510)" to="(3650,530)"/>
    <wire from="(3650,530)" to="(3690,530)"/>
    <wire from="(3650,550)" to="(3650,1380)"/>
    <wire from="(3660,540)" to="(3660,610)"/>
    <wire from="(3660,540)" to="(3690,540)"/>
    <wire from="(3670,550)" to="(3670,640)"/>
    <wire from="(3670,550)" to="(3690,550)"/>
    <wire from="(3680,580)" to="(3680,1100)"/>
    <wire from="(3680,580)" to="(3690,580)"/>
    <wire from="(3690,600)" to="(3690,1400)"/>
    <wire from="(3710,560)" to="(3710,570)"/>
    <wire from="(3730,540)" to="(3740,540)"/>
    <wire from="(3740,540)" to="(3740,1410)"/>
    <wire from="(420,600)" to="(430,600)"/>
    <wire from="(430,290)" to="(430,560)"/>
    <wire from="(430,290)" to="(500,290)"/>
    <wire from="(430,560)" to="(430,600)"/>
    <wire from="(430,560)" to="(760,560)"/>
    <wire from="(470,600)" to="(480,600)"/>
    <wire from="(70,150)" to="(1550,150)"/>
    <wire from="(70,150)" to="(70,370)"/>
    <wire from="(70,870)" to="(100,870)"/>
    <wire from="(720,290)" to="(730,290)"/>
    <wire from="(720,650)" to="(730,650)"/>
    <wire from="(730,210)" to="(730,290)"/>
    <wire from="(730,290)" to="(1530,290)"/>
    <wire from="(730,290)" to="(730,580)"/>
    <wire from="(730,580)" to="(760,580)"/>
    <wire from="(730,620)" to="(730,650)"/>
    <wire from="(730,620)" to="(760,620)"/>
    <wire from="(750,1300)" to="(1170,1300)"/>
    <wire from="(750,520)" to="(1640,520)"/>
    <wire from="(750,520)" to="(750,540)"/>
    <wire from="(750,540)" to="(760,540)"/>
    <wire from="(750,600)" to="(750,1300)"/>
    <wire from="(750,600)" to="(760,600)"/>
    <wire from="(760,1160)" to="(1170,1160)"/>
    <wire from="(760,1160)" to="(760,1400)"/>
    <wire from="(760,1400)" to="(940,1400)"/>
    <wire from="(770,1150)" to="(1160,1150)"/>
    <wire from="(770,1150)" to="(770,1380)"/>
    <wire from="(770,1380)" to="(940,1380)"/>
    <wire from="(790,1280)" to="(1990,1280)"/>
    <wire from="(790,1280)" to="(790,1360)"/>
    <wire from="(790,1360)" to="(940,1360)"/>
    <wire from="(80,400)" to="(80,640)"/>
    <wire from="(80,640)" to="(200,640)"/>
    <wire from="(830,1320)" to="(830,1460)"/>
    <wire from="(830,1320)" to="(940,1320)"/>
    <wire from="(830,1460)" to="(1240,1460)"/>
    <wire from="(860,1250)" to="(1890,1250)"/>
    <wire from="(860,1250)" to="(860,1340)"/>
    <wire from="(860,1340)" to="(940,1340)"/>
    <wire from="(90,210)" to="(730,210)"/>
    <wire from="(90,210)" to="(90,370)"/>
    <wire from="(90,620)" to="(130,620)"/>
    <wire from="(90,620)" to="(90,890)"/>
    <wire from="(90,890)" to="(240,890)"/>
    <wire from="(980,540)" to="(1660,540)"/>
    <wire from="(980,560)" to="(990,560)"/>
    <wire from="(980,580)" to="(1000,580)"/>
    <wire from="(990,560)" to="(990,890)"/>
    <wire from="(990,890)" to="(1620,890)"/>
  </circuit>


  <vhdl name="ALU">library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.ALL;
USE IEEE.std_logic_unsigned.ALL;

entity ALU is
    port(
    A, B      : in std_logic_vector(31 downto 0);  -- Entradas A e B de 32 bits
    control   : in std_logic_vector(3 downto 0);   -- Entrada de controle de 4 bits
    result    : out std_logic_vector(31 downto 0); -- Saída de resultado de 32 bits
    zero      : out std_logic);                    -- Saída para sinalizar se o resultado é zero
end ALU;

architecture TypeArchitecture of ALU is

signal zero_out   : std_logic_vector(32 downto 0); -- Vetor para verificação de resultado zero
signal result_out : std_logic_vector(31 downto 0); -- Vetor para armazenar o resultado da operação

begin
	
    result_out &lt;= (A + B) when control = "0010" else                  -- Soma
    			   (A - B) when control = "0110" else                  -- Subtração
    			   (A XOR B) when control = "0101" else                -- XOR (ou exclusivo)
    			   (A OR B) when control = "0001" else                 -- OR (ou)
    			   (A AND B) when control = "0000" else                -- AND (e)
    			   (std_logic_vector(shift_left(unsigned(A), to_integer(unsigned(B))))) when control = "0011" else   -- Shift Left (deslocamento à esquerda)
    			   (std_logic_vector(shift_right(unsigned(A), to_integer(unsigned(B))))) when control = "0111";    -- Shift Right (deslocamento à direita)
        			
    result &lt;= result_out;                          -- Atribui o valor do resultado à saída result
    zero_out(0) &lt;= '0';                            -- Inicializa o primeiro bit de zero_out como '0'
    G2: for I in 1 to 32 generate
            zero_out(I) &lt;= zero_out(I - 1) or result_out(I - 1);  -- Verificação de resultado zero bit a bit
    end generate;
    zero &lt;= not zero_out(32);                      -- Sinaliza se o resultado é zero (se zero_out(32) for '0', zero é '1', caso contrário, zero é '0')
end TypeArchitecture;
</vhdl>


  <vhdl name="ALU_Control">library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ALU_Control is
    port(
        Functs    : IN std_logic_vector(3 downto 0);    -- Entrada de códigos de função da ALU (4 bits)
        AluOp   : IN std_logic_vector(1 downto 0);      -- Entrada de códigos de operação da ALU (2 bits)
        Control : OUT std_logic_vector(3 downto 0)      -- Saída do controle da ALU (4 bits)
        );
end ALU_Control;

architecture TypeArchitecture of ALU_Control is
begin

	control &lt;= "0010" when AluOp = "00" else -- Se AluOp for "00", Control recebe "0010" (Operação: Soma)
			 "0110" when AluOp = "01" else -- Se AluOp for "01", Control recebe "0110" (Operação: Branch)
			 "0010" when Functs = "0000" else -- Se Functs for "0000", Control recebe "0010" (Operação: Adição)
			 "0110" when Functs = "1000" else -- Se Functs for "1000", Control recebe "0110" (Operação: Subtração)
			 "0011" when Functs = "0001" else -- Se Functs for "0001", Control recebe "0011" (Operação: Shift Left)
			 "0101" when Functs = "0100" else -- Se Functs for "0100", Control recebe "0101" (Operação: XOR)
			 "0111" when Functs = "0101" else -- Se Functs for "0101", Control recebe "0111" (Operação: Shift Right)
			 "0001" when Functs = "0110" else -- Se Functs for "0110", Control recebe "0001" (Operação: OR)
			 "0000" when Functs = "0111"; -- Se Functs for "0111", Control recebe "0000" (Operação: AND)
	 
end TypeArchitecture;
</vhdl>
  <vhdl name="Control_Unit">library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Control_Unit is
    port(
        opcode                     : IN  std_logic_vector(6 downto 0);  -- Entrada do código de operação (7 bits)
        AluSrc, blockA, RegWrite   : OUT std_logic;                      -- Saída de sinais de controle individuais (1 bit cada)
        MemRead, MemWrite, Branch  : OUT std_logic;                      -- Saída de sinais de controle individuais (1 bit cada)
        BranchNotEq, BrIncond      : OUT std_logic;                      -- Saída de sinais de controle individuais (1 bit cada)
        regToPC                    : OUT std_logic;                      -- Saída de sinal de controle (1 bit)
        AluOp, regSrc              : OUT std_logic_vector(1 downto 0)    -- Saída de códigos de operação da ALU e seleção de registradores (2 bits cada)
        );
end Control_Unit;

architecture TypeArchitecture of Control_Unit is
begin
    -- Processo que verifica o opcode e define os sinais de controle correspondentes
    process(opcode)
    begin
        IF (opcode = "0110011") THEN -- R-Type sem imediato (add, sub, and, or, xor, slt)
            AluSrc      &lt;= '0';  -- Seleção de fonte para a ALU (0: A_i, 1: Immediato)
            blockA      &lt;= '0';  -- Seleção de origem do registrador A (0: rs1, 1: zero)
            RegWrite    &lt;= '1';  -- Habilita escrita no registrador destino
            MemRead     &lt;= '0';  -- Habilita leitura de memória
            MemWrite    &lt;= '0';  -- Habilita escrita na memória
            Branch      &lt;= '0';  -- Habilita desvio condicional
            AluOp       &lt;= "10"; -- Código de operação da ALU para R-Type (00: and, 01: or, 10: add, 11: sub)
            regSrc      &lt;= "00"; -- Seleção de registradores para R-Type (00: rs1, 01: rs2, 10: rd, 11: zero)
            BranchNotEq &lt;= '0';  -- Habilita desvio condicional se as entradas forem diferentes
            BrIncond    &lt;= '0';  -- Habilita desvio incondicional
            regToPC     &lt;= '0';  -- Seleção de registrador para atualizar o PC (0: PC+4, 1: rd)
        END IF;

        IF (opcode = "0010011") THEN -- I-Type (addi, andi, ori, xori, slti)
            AluSrc      &lt;= '1';  -- Seleção de fonte para a ALU (0: A_i, 1: Immediato)
            blockA      &lt;= '0';  -- Seleção de origem do registrador A (0: rs1, 1: zero)
            RegWrite    &lt;= '1';  -- Habilita escrita no registrador destino
            MemRead     &lt;= '0';  -- Habilita leitura de memória
            MemWrite    &lt;= '0';  -- Habilita escrita na memória
            Branch      &lt;= '0';  -- Habilita desvio condicional
            AluOp       &lt;= "11"; -- Código de operação da ALU para I-Type (00: andi, 01: ori, 10: addi, 11: slti)
            regSrc      &lt;= "00"; -- Seleção de registradores para I-Type (00: rs1, 01: rd, 10: zero)
            BranchNotEq &lt;= '0';  -- Habilita desvio condicional se as entradas forem diferentes
            BrIncond    &lt;= '0';  -- Habilita desvio incondicional
            regToPC     &lt;= '0';  -- Seleção de registrador para atualizar o PC (0: PC+4, 1: rd)
        END IF;

        IF (opcode = "0100011") THEN -- S-Type (sw)
            AluSrc      &lt;= '1';  -- Seleção de fonte para a ALU (0: A_i, 1: Immediato)
            blockA      &lt;= '0';  -- Seleção de origem do registrador A (0: rs1, 1: zero)
            RegWrite    &lt;= '0';  -- Habilita escrita no registrador destino
            MemRead     &lt;= '0';  -- Habilita leitura de memória
            MemWrite    &lt;= '1';  -- Habilita escrita na memória
            Branch      &lt;= '0';  -- Habilita desvio condicional
            AluOp       &lt;= "00"; -- Código de operação da ALU para S-Type (00: add)
            regSrc      &lt;= "00"; -- Seleção de registradores para S-Type (00: rs1, 01: zero)
            BranchNotEq &lt;= '0';  -- Habilita desvio condicional se as entradas forem diferentes
            BrIncond    &lt;= '0';  -- Habilita desvio incondicional
            regToPC     &lt;= '0';  -- Seleção de registrador para atualizar o PC (0: PC+4, 1: rd)
        END IF;

        IF (opcode = "1100111") THEN -- SB-Type (beq)
            AluSrc      &lt;= '0';  -- Seleção de fonte para a ALU (0: A_i, 1: Immediato)
            blockA      &lt;= '0';  -- Seleção de origem do registrador A (0: rs1, 1: zero)
            RegWrite    &lt;= '0';  -- Habilita escrita no registrador destino
            MemRead     &lt;= '0';  -- Habilita leitura de memória
            MemWrite    &lt;= '0';  -- Habilita escrita na memória
            Branch      &lt;= '1';  -- Habilita desvio condicional
            AluOp       &lt;= "01"; -- Código de operação da ALU para SB-Type (01: sub)
            regSrc      &lt;= "00"; -- Seleção de registradores para SB-Type (00: rs1, 01: rs2)
            BranchNotEq &lt;= '0';  -- Habilita desvio condicional se as entradas forem diferentes
            BrIncond    &lt;= '0';  -- Habilita desvio incondicional
            regToPC     &lt;= '0';  -- Seleção de registrador para atualizar o PC (0: PC+4, 1: rd)
        END IF;

        IF (opcode = "1100011") THEN -- SB-Type (bne)
            AluSrc      &lt;=
</vhdl>
  <vhdl name="ImmGen">library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity ImmGen is
    Port( 
        inst: in std_logic_vector(31 downto 0);  -- Entrada da instrução (32 bits)
        imm: out std_logic_vector(31 downto 0)  -- Saída do valor imediato gerado (32 bits)
        );
end ImmGen;

architecture Behavioral of ImmGen is
    signal opcode       : std_logic_vector(6 downto 0);  -- Sinal para armazenar o campo opcode da instrução (7 bits)
    signal imm_interno  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";  -- Valor imediato interno inicializado com zero

begin

    opcode &lt;= inst(6 downto 0);  -- Extrai o campo opcode da instrução

    process(opcode)
    begin
        if (opcode = "0010011" or opcode = "1100110") then  -- Tipo I (load-immediate, jump-register)
            imm_interno(11 downto 0)  &lt;= inst(31 downto 20);  -- Extrai o imediato de 11 bits
            imm_interno(31 downto 12) &lt;= (others =&gt; inst(31));  -- Sinal extendido para os bits mais significativos
        elsif (opcode = "1110111" or opcode = "0110111") then  -- Tipo U (lui, auipc)
            imm_interno(31 downto 12) &lt;= inst(31 downto 12);  -- Extrai o imediato de 20 bits
        elsif (opcode = "0100011") then  -- Tipo S (store)
            imm_interno(11 downto 5)  &lt;= inst(31 downto 25);  -- Extrai o imediato de 7 bits (5-11)
            imm_interno(4 downto 0)   &lt;= inst(11 downto 7);   -- Extrai o imediato de 5 bits (0-4)
            imm_interno(31 downto 12) &lt;= (others =&gt; inst(31));  -- Sinal extendido para os bits mais significativos
        elsif (opcode = "1100111" or opcode = "1100011") then  -- Tipo SB (branch)
            imm_interno(12)           &lt;= inst(31);          -- Extrai o bit de imediato (12)
            imm_interno(11)           &lt;= inst(7);           -- Extrai o bit de imediato (11)
            imm_interno(10 downto 5)  &lt;= inst(30 downto 25);  -- Extrai o imediato de 6 bits (5-10)
            imm_interno(4 downto 1)   &lt;= inst(11 downto 8);   -- Extrai o imediato de 4 bits (1-4)
            imm_interno(31 downto 13) &lt;= (others =&gt; inst(31));  -- Sinal extendido para os bits mais significativos
        elsif (opcode = "1101111") then  -- Tipo UJ (jump)
            imm_interno(20)           &lt;= inst(31);          -- Extrai o bit de imediato (20)
            imm_interno(19 downto 12) &lt;= inst(19 downto 12);  -- Extrai o imediato de 8 bits (12-19)
            imm_interno(11)           &lt;= inst(20);          -- Extrai o bit de imediato (11)
            imm_interno(10 downto 1)  &lt;= inst(30 downto 21);  -- Extrai o imediato de 10 bits (1-10)
        end if;
    end process;

    imm &lt;= imm_interno;  -- Define a saída como o valor imediato gerado

end Behavioral;
</vhdl>
  <vhdl name="PC2">LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY PC2 IS
  PORT (
  ------------------------------------------------------------------------------
  --Insert input ports below
    clk      : IN  std_logic;                    -- Entrada do sinal de clock
    reset    : IN  std_logic;                    -- Entrada do sinal de reset
    pc_in    : IN  std_logic_vector(31 DOWNTO 0); -- Entrada do valor atual do PC (contador de programa)
    writeEnableL   : IN std_logic;               -- Entrada do sinal de habilitação de escrita no PC
  ------------------------------------------------------------------------------
  --Insert output ports below
    pc_out   : OUT std_logic_vector(31 DOWNTO 0)  -- Saída do valor atualizado do PC (contador de programa)
    );
END PC2;

--------------------------------------------------------------------------------
--Complete your VHDL description below
--------------------------------------------------------------------------------

ARCHITECTURE TypeArchitecture OF PC2 IS

BEGIN

	
	PROCESS (clk, reset, writeEnableL)
	BEGIN
		IF (rising_edge(clk)) THEN                      -- Detecta a borda de subida do sinal de clock
			if (pc_in = "UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU") then   -- Verifica se o valor atual do PC é desconhecido (não inicializado)
				pc_out &lt;= (others =&gt; '0');               -- Se for desconhecido, zera o valor do PC
			elsif (writeEnableL = '0') then              -- Verifica se o sinal de habilitação de escrita está desabilitado
				pc_out &lt;= pc_in;                         -- Se estiver desabilitado, o PC mantém o valor atual (não ocorre atualização)
			end if;
		END IF;
		IF (reset = '1') THEN                           -- Detecta a ocorrência de um reset (sinal de reset em nível alto)
			pc_out &lt;= (others =&gt; '0');                   -- Nesse caso, zera o valor do PC
		END IF;
	END PROCESS;

END TypeArchitecture;
</vhdl>
  <vhdl name="somador">LIBRARY ieee;
USE ieee.std_logic_1164.all;

USE IEEE.std_logic_unsigned.ALL; -- Pacote para operações aritméticas com std_logic_vector

ENTITY somador IS
  PORT (
  ------------------------------------------------------------------------------
    A, B        : IN  std_logic_vector(31 DOWNTO 0); -- Vetor de entrada exemplo A e B de 32 bits
  ------------------------------------------------------------------------------
    Z           : OUT std_logic_vector(31 DOWNTO 0)  -- Vetor de saída exemplo Z de 32 bits
    );
END somador;

ARCHITECTURE TypeArchitecture OF somador IS

BEGIN

Z &lt;= A + B; -- Saída Z é a soma dos vetores de entrada A e B

END TypeArchitecture;
</vhdl>
  <vhdl name="register_file">library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity register_file is
  port(
    outA        : out std_logic_vector(31 downto 0);    -- Saída A do registrador
    outB        : out std_logic_vector(31 downto 0);    -- Saída B do registrador
    input       : in  std_logic_vector(31 downto 0);    -- Entrada de dado para escrita no registrador
    regSelManual: in  std_logic_vector(4 downto 0);     -- Seleção manual de um registrador de saída
    outRegManual: out std_logic_vector(31 downto 0);    -- Saída do registrador selecionado manualmente
    writeEnable : in  std_logic;                        -- Sinal de habilitação de escrita no registrador
    regASel     : in  std_logic_vector(4 downto 0);     -- Seleção do registrador A para leitura
    regBSel     : in  std_logic_vector(4 downto 0);     -- Seleção do registrador B para leitura
    writeRegSel : in  std_logic_vector(4 downto 0);     -- Seleção do registrador para escrita
    clk         : in  std_logic                        -- Sinal de clock
    );
end register_file;

architecture TypeArchitecture of register_file is
  type registerFile is array(0 to 31) of std_logic_vector(31 downto 0);
  signal registers : registerFile := 
   -- Valores iniciais dos registradores
   -- Os primeiros 32 registradores têm os valores pré-definidos como "00000000000000000000000000010000", "00000000000000000000000000000001", etc.
   -- Até o último registrador "00000000000000000000000000000000"
   ("00000000000000000000000000010000","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000");

begin
  regFile : process (clk) is
  begin
    if rising_edge(clk) then
      -- Read A and B before bypass
      -- Leitura dos registradores A e B antes do bypass
      if (registers(to_integer(unsigned(regASel))) = "UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU") THEN
      	outA &lt;= (others =&gt; '0');  -- Se o valor for "UUUU..." (indeterminado), a saída A será "0000..."
      ELSE 
      	outA &lt;= registers(to_integer(unsigned(regASel)));  -- Caso contrário, a saída A será o valor do registrador selecionado
      END IF;
      IF (registers(to_integer(unsigned(regBSel))) = "UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU") THEN
      	outB &lt;= (others =&gt; '0');  -- Se o valor for "UUUU..." (indeterminado), a saída B será "0000..."
      ELSE
      	outB &lt;= registers(to_integer(unsigned(regBSel)));  -- Caso contrário, a saída B será o valor do registrador selecionado
      END IF;
      -- Write and bypass
      -- Escrita e bypass
      if writeEnable = '1' then
        registers(to_integer(unsigned(writeRegSel))) &lt;= input;  -- Escreve o valor da entrada no registrador selecionado
        if regASel = writeRegSel then  -- Bypass para leitura A
          outA &lt;= input;  -- Se o registrador A é o mesmo selecionado para escrita, a saída A recebe o valor da entrada
        end if;
        if regBSel = writeRegSel then  -- Bypass para leitura B
          outB &lt;= input;  -- Se o registrador B é o mesmo selecionado para escrita, a saída B recebe o valor da entrada
        end if;
      end if;
    end if;
  end process;

  -- seleção manual
  -- O valor de saída outRegManual recebe o valor do registrador selecionado manualmente (regSelManual)
  outRegManual &lt;= registers(to_integer(unsigned(regSelManual)));
  
end TypeArchitecture;
</vhdl>
  <vhdl name="IFID">LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY IFID IS
  PORT (
    clk         : IN  std_logic;                    -- Entrada do sinal de clock
    pcIn        : IN  std_logic_vector(31 DOWNTO 0); -- Entrada do valor atual do PC (contador de programa)
    pcPl4In	 : IN  std_logic_vector(31 downto 0); -- Entrada do valor do PC mais 4 (próxima instrução)
    writeEnableL   : IN std_logic;                 -- Entrada do sinal de habilitação de escrita no IFID
    instIn      : IN  std_logic_vector(31 DOWNTO 0); -- Entrada da instrução atual buscada na memória de instruções
    pcOut       : OUT std_logic_vector(31 DOWNTO 0); -- Saída do valor atual do PC (contador de programa)
    pcPl4Out	 : OUT std_logic_vector(31 downto 0); -- Saída do valor do PC mais 4 (próxima instrução)
    instOut     : OUT std_logic_vector(31 DOWNTO 0)  -- Saída da instrução atual buscada na memória de instruções
    );
END IFID;


ARCHITECTURE TypeArchitecture OF IFID IS

SIGNAL IDIF : std_logic_vector(95 DOWNTO 0);  -- Registrador de 96 bits para armazenar os valores do IFID

BEGIN


	
	PROCESS (clk, writeEnableL)
	BEGIN
		IF (rising_edge(clk)) THEN                   -- Detecta a borda de subida do sinal de clock
			if (writeEnableL = '0') then             -- Verifica se o sinal de habilitação de escrita está desabilitado
				IDIF(31 DOWNTO 0) &lt;= instIn;         -- Se estiver desabilitado, armazena a instrução atual no IFID
				IDIF(63 DOWNTO 32) &lt;= pcIn;          -- Armazena o valor atual do PC
				IDIF(95 downto 64) &lt;= pcPl4In;       -- Armazena o valor do PC mais 4 (próxima instrução)
			end if;
		END IF;
		IF (falling_edge(clk)) THEN                 -- Detecta a borda de descida do sinal de clock
			pcOut &lt;= IDIF(63 DOWNTO 32);           -- Na borda de descida, coloca na saída o valor do PC atual
			instOut &lt;= IDIF(31 DOWNTO 0);          -- Coloca na saída a instrução armazenada no IFID
			pcPl4Out &lt;= IDIF(95 downto 64);        -- Coloca na saída o valor do PC mais 4
		END IF;
	END PROCESS;

	
END TypeArchitecture;
</vhdl>
  <vhdl name="IDEX">LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY IDEX IS
  PORT (
    clk            : IN  std_logic;                    -- Entrada do sinal de clock
    pcIn           : IN  std_logic_vector(31 DOWNTO 0); -- Entrada do valor atual do PC (contador de programa)
    read1In        : IN  std_logic_vector(31 DOWNTO 0); -- Entrada do valor lido do registrador 1
    read2In        : IN  std_logic_vector(31 DOWNTO 0); -- Entrada do valor lido do registrador 2
    immGenIn       : in  std_logic_vector(31 DOWNTO 0); -- Entrada do valor gerado pela unidade ImmGen
    aluControlin   : IN  std_logic_vector(3 downto 0);  -- Entrada do controle da ALU
    wbAddIn        : IN  std_logic_vector(4 downto 0);  -- Entrada do endereço do registrador de destino para escrita
    WBin		    : IN  std_logic_vector(2 downto 0);  -- Entrada da fonte de escrita no registrador de destino
    Min 		    : IN  std_logic_vector(5 downto 0);  -- Entrada do sinal de controle de escrita na memória de dados
    EXin    	    : IN  std_logic_vector(3 downto 0);  -- Entrada do sinal de controle de execução
    pcPl4In	    : IN  std_logic_vector(31 downto 0); -- Entrada do valor do PC mais 4 (próxima instrução)
    rs1In		    : IN  std_logic_vector(4 downto 0);  -- Entrada do endereço do registrador 1
    rs2In		    : IN  std_logic_vector(4 downto 0);  -- Entrada do endereço do registrador 2
                        
    pcOut          : OUT std_logic_vector(31 DOWNTO 0); -- Saída do valor atual do PC (contador de programa)
    read1Out	    : OUT std_logic_vector(31 DOWNTO 0); -- Saída do valor lido do registrador 1
    read2Out       : OUT std_logic_vector(31 DOWNTO 0); -- Saída do valor lido do registrador 2
    immGenOut      : OUT std_logic_vector(31 DOWNTO 0); -- Saída do valor gerado pela unidade ImmGen
    aluControlout  : OUT std_logic_vector(3 downto 0);  -- Saída do controle da ALU
    wbAddOut       : OUT std_logic_vector(4 downto 0);  -- Saída do endereço do registrador de destino para escrita
    WBout		    : OUT std_logic_vector(2 downto 0);  -- Saída da fonte de escrita no registrador de destino
    Mout 		    : OUT std_logic_vector(5 downto 0);  -- Saída do sinal de controle de escrita na memória de dados
    EXout    	    : OUT std_logic_vector(3 downto 0);  -- Saída do sinal de controle de execução
    pcPl4Out	    : OUT std_logic_vector(31 downto 0); -- Saída do valor do PC mais 4 (próxima instrução)
    rs1Out	    : OUT std_logic_vector(4 downto 0);  -- Saída do endereço do registrador 1
    rs2Out	    : OUT std_logic_vector(4 downto 0)   -- Saída do endereço do registrador 2
    );
END IDEX;


ARCHITECTURE TypeArchitecture OF IDEX IS

SIGNAL idex_s : std_logic_vector(191 DOWNTO 0);  -- Registrador de 192 bits para armazenar os valores do IDEX

BEGIN

	PROCESS (clk)
	BEGIN
		IF (rising_edge(clk)) THEN                   -- Detecta a borda de subida do sinal de clock
			idex_s(31 DOWNTO 0)    &lt;= pcIn;          -- Armazena o valor atual do PC
			idex_s(63 DOWNTO 32)   &lt;= read1In;       -- Armazena o valor lido do registrador 1
			idex_s(95 DOWNTO 64)   &lt;= read2In;       -- Armazena o valor lido do registrador 2
			idex_s(127 DOWNTO 96)  &lt;= immGenIn;      -- Armazena o valor gerado pela unidade ImmGen
			idex_s(131 DOWNTO 128) &lt;= aluControlin;  -- Armazena o controle da ALU
			idex_s(136 DOWNTO 132) &lt;= wbAddIn;       -- Armazena o endereço do registrador de destino para escrita
			idex_s(139 downto 137) &lt;= WBin;          -- Armazena a fonte de escrita no registrador de destino
			idex_s(145 downto 140) &lt;= Min;           -- Armazena o sinal de controle de escrita na memória de dados
			idex_s(149 downto 146) &lt;= EXin;          -- Armazena o sinal de controle de execução
			idex_s(181 downto 150) &lt;= pcPl4In;       -- Armazena o valor do PC mais 4 (próxima instrução)
			idex_s(186 downto 182) &lt;= rs1In;         -- Armazena o endereço do registrador 1
			idex_s(191 downto 187) &lt;= rs2In;         -- Armazena o endereço do registrador 2
		END IF;
		IF (falling_edge(clk)) THEN                 -- Detecta a borda de descida do sinal de clock
			pcOut    &lt;= idex_s(31 DOWNTO 0);        -- Na borda de descida, coloca na saída o valor do PC atual
			read1Out  &lt;= idex_s(63 DOWNTO 32);      -- Coloca na saída o valor lido do registrador 1
			read2Out  &lt;= idex_s(95 DOWNTO 64);      -- Coloca na saída o valor lido do registrador 2
			immGenOut &lt;= idex_s(127 DOWNTO 96);     -- Coloca na saída
			aluControlout &lt;= idex_s(131 DOWNTO 128);
			wbAddOut &lt;= idex_s(136 DOWNTO 132);
			WBout &lt;= idex_s(139 downto 137);
			Mout &lt;= idex_s(145 downto 140);
			EXout &lt;= idex_s(149 downto 146);
			pcPl4Out &lt;= idex_s(181 downto 150);
			rs1Out &lt;= idex_s(186 downto 182);
			rs2Out &lt;= idex_s(191 downto 187);
		END IF;
	END PROCESS;

	
END TypeArchitecture;
</vhdl>
  <vhdl name="EXMEM">LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY EXMEM IS
  PORT (
    clk            : IN  std_logic;                    -- Entrada do sinal de clock
    sumIn           : IN  std_logic_vector(31 DOWNTO 0); -- Entrada do resultado da ALU
    zeroIn        : IN  std_logic;                    -- Entrada do sinal de zero da ALU
    aluIn        : IN  std_logic_vector(31 DOWNTO 0);  -- Entrada da operação da ALU
    read2In       : IN  std_logic_vector(31 DOWNTO 0);  -- Entrada do valor lido do registrador 2
    wbAddIn        : IN  std_logic_vector(4 downto 0);  -- Entrada do endereço do registrador de destino para escrita
    WBin		    : IN  std_logic_vector(2 downto 0);  -- Entrada da fonte de escrita no registrador de destino
    Min 		    : IN  std_logic_vector(5 downto 0);  -- Entrada do sinal de controle de escrita na memória de dados
    pcPl4In	    : IN std_logic_vector(31 downto 0);  -- Entrada do valor do PC mais 4 (próxima instrução)
    
    pcOut         : OUT std_logic_vector(31 DOWNTO 0); -- Saída do valor atual do PC (contador de programa)
    zeroOut	    : OUT std_logic;                    -- Saída do sinal de zero da ALU
    aluOut       : OUT std_logic_vector(31 DOWNTO 0);  -- Saída do resultado da ALU
    read2Out      : OUT std_logic_vector(31 DOWNTO 0); -- Saída do valor lido do registrador 2
    wbAddOut       : OUT std_logic_vector(4 downto 0);  -- Saída do endereço do registrador de destino para escrita
    WBout		    : OUT std_logic_vector(2 downto 0);  -- Saída da fonte de escrita no registrador de destino
    Mout 		    : OUT std_logic_vector(5 downto 0);  -- Saída do sinal de controle de escrita na memória de dados
    pcPl4Out	    : OUT std_logic_vector(31 downto 0)  -- Saída do valor do PC mais 4 (próxima instrução)
    );
END EXMEM;


ARCHITECTURE TypeArchitecture OF EXMEM IS

SIGNAL exmem_s : std_logic_vector(142 DOWNTO 0);  -- Registrador de 143 bits para armazenar os valores do EXMEM

BEGIN

	PROCESS (clk)
	BEGIN
		IF (rising_edge(clk)) THEN                    -- Detecta a borda de subida do sinal de clock
			exmem_s(31 DOWNTO 0)   &lt;= sumIn;          -- Armazena o resultado da ALU
			exmem_s(32)  &lt;= zeroIn;                   -- Armazena o sinal de zero da ALU
			exmem_s(64 DOWNTO 33)  &lt;= aluIn;          -- Armazena a operação da ALU
			exmem_s(96 DOWNTO 65) &lt;= read2In;         -- Armazena o valor lido do registrador 2
			exmem_s(101 DOWNTO 97) &lt;= wbAddIn;        -- Armazena o endereço do registrador de destino para escrita
			exmem_s(104 DOWNTO 102) &lt;= WBin;          -- Armazena a fonte de escrita no registrador de destino
			exmem_s(110 DOWNTO 105) &lt;= Min;           -- Armazena o sinal de controle de escrita na memória de dados
			exmem_s(142 downto 111) &lt;= pcPl4In;       -- Armazena o valor do PC mais 4 (próxima instrução)
		END IF;
		IF (falling_edge(clk)) THEN                  -- Detecta a borda de descida do sinal de clock
			pcOut    &lt;=  exmem_s(31 DOWNTO 0);       -- Na borda de descida, coloca na saída o valor do PC atual
			zeroOut  &lt;=  exmem_s(32);                -- Coloca na saída o sinal de zero da ALU
			aluOut   &lt;=  exmem_s(64 DOWNTO 33);       -- Coloca na saída o resultado da ALU
			read2Out &lt;=  exmem_s(96 DOWNTO 65);       -- Coloca na saída o valor lido do registrador 2
			wbAddOut &lt;=  exmem_s(101 DOWNTO 97);      -- Coloca na saída o endereço do registrador de destino para escrita
			WBout    &lt;=  exmem_s(104 DOWNTO 102);     -- Coloca na saída a fonte de escrita no registrador de destino
			Mout     &lt;=  exmem_s(110 DOWNTO 105);     -- Coloca na saída o sinal de controle de escrita na memória de dados
			pcPl4Out &lt;=  exmem_s(142 downto 111);     -- Coloca na saída o valor do PC mais 4 (próxima instrução)
		END IF;
	END PROCESS;

	
END TypeArchitecture;
</vhdl>
  <vhdl name="MEMWB">LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY MEMWB IS
  PORT (
    clk            : IN  std_logic;                    -- Entrada do sinal de clock
    readIn         : IN  std_logic_vector(31 DOWNTO 0); -- Entrada do valor lido da memória ou resultado da ALU
    aluIn          : IN  std_logic_vector(31 DOWNTO 0); -- Entrada do resultado da operação da ALU
    wbAddIn        : IN  std_logic_vector(4 downto 0);  -- Entrada do endereço do registrador de destino para escrita
    WBin		    : IN  std_logic_vector(2 downto 0);  -- Entrada da fonte de escrita no registrador de destino
    pcPl4In	    : IN std_logic_vector(31 downto 0); -- Entrada do valor do PC mais 4 (próxima instrução)
    pcPlIIn	    : IN std_logic_vector(31 downto 0); -- Entrada do valor do PC mais I (endereço de retorno para chamadas de função)
                        
    readOut        : OUT std_logic_vector(31 DOWNTO 0); -- Saída do valor lido da memória ou resultado da ALU
    aluOut	        : OUT std_logic_vector(31 DOWNTO 0); -- Saída do resultado da operação da ALU
    wbAddOut       : OUT std_logic_vector(4 downto 0);  -- Saída do endereço do registrador de destino para escrita
    WBout		    : OUT std_logic_vector(2 downto 0);  -- Saída da fonte de escrita no registrador de destino
    pcPl4Out       : OUT std_logic_vector(31 downto 0); -- Saída do valor do PC mais 4 (próxima instrução)
    pcPlIOut	    : OUT std_logic_vector(31 downto 0)  -- Saída do valor do PC mais I (endereço de retorno para chamadas de função)
    );
END MEMWB;

ARCHITECTURE TypeArchitecture OF MEMWB IS

SIGNAL memwb_s : std_logic_vector(135 DOWNTO 0);  -- Registrador de 136 bits para armazenar os valores do MEMWB

BEGIN

	PROCESS (clk)
	BEGIN
		IF (rising_edge(clk)) THEN                       -- Detecta a borda de subida do sinal de clock
			memwb_s(31 DOWNTO 0)   &lt;= readIn;            -- Armazena o valor lido da memória ou resultado da ALU
			memwb_s(63 DOWNTO 32)  &lt;= aluIn;             -- Armazena o resultado da operação da ALU
			memwb_s(68 DOWNTO 64)  &lt;= wbAddIn;           -- Armazena o endereço do registrador de destino para escrita
			memwb_s(71 DOWNTO 69)  &lt;= WBin;              -- Armazena a fonte de escrita no registrador de destino
			memwb_s(103 downto 72) &lt;= pcPl4In;           -- Armazena o valor do PC mais 4 (próxima instrução)
			memwb_s(135 downto 104) &lt;= pcPlIIn;          -- Armazena o valor do PC mais I (endereço de retorno para chamadas de função)
			
		END IF;
		IF (falling_edge(clk)) THEN                      -- Detecta a borda de descida do sinal de clock
			readOut    &lt;=  memwb_s(31 DOWNTO 0);         -- Na borda de descida, coloca na saída o valor lido da memória ou resultado da ALU
			aluOut     &lt;=  memwb_s(63 DOWNTO 32);        -- Coloca na saída o resultado da operação da ALU
			wbAddOut   &lt;=  memwb_s(68 DOWNTO 64);        -- Coloca na saída o endereço do registrador de destino para escrita
			WBout      &lt;=  memwb_s(71 DOWNTO 69);        -- Coloca na saída a fonte de escrita no registrador de destino
			pcPl4Out   &lt;=  memwb_s(103 downto 72);       -- Coloca na saída o valor do PC mais 4 (próxima instrução)
			pcPlIOut   &lt;=  memwb_s(135 downto 104);      -- Coloca na saída o valor do PC mais I (endereço de retorno para chamadas de função)
		END IF;
	END PROCESS;

	
END TypeArchitecture;
</vhdl>
  <vhdl name="Harzard">library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Harzard is 
	port( 
        clk 		   : IN std_logic;                          -- Entrada do sinal de clock
        MemReadEX 	   : IN std_logic;                          -- Sinal indicando leitura na memória (saída do estágio EX do pipeline)
        RDEX, RSrc1, RSrc2 : IN std_logic_vector(4 downto 0);  -- Registradores de destino e fontes da instrução (saídas do estágio EX do pipeline)
        stall		   : OUT std_logic                         -- Saída que indica se um "stall" (atraso) deve ser aplicado
	);
end Harzard;

architecture TypeArchitecture of Harzard is
	signal stall_interno : std_logic := '0';  -- Sinal interno que armazena o valor do stall

begin
	process(clk)
    begin
        if ((MemReadEX = '1') and ((RDEX = RSrc1) or (RDEX = RSrc2))) then
            stall_interno &lt;='1';  -- Se houver uma leitura na memória (MemReadEX = '1') e o resultado da EX estiver em RSrc1 ou RSrc2, aplica um stall
        end if;
    end process;
    stall &lt;= stall_interno;  -- Atribui o valor do sinal interno stall_interno à saída stall
end TypeArchitecture;
</vhdl>
  <vhdl name="Forward">library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Forward is 
	port( 
	     clk					: IN std_logic;                      -- Entrada do sinal de clock
	     regWriteWB, regWriteMEM 	: IN std_logic;                      -- Sinais de escrita no registrador (saídas de MEM/WB e WB do pipeline)
	     RSrc1, RSrc2			: IN std_logic_vector(4 downto 0);   -- Registradores fonte da instrução (saídas de ID/EX do pipeline)
	     RDWB, RDMEM			: IN std_logic_vector(4 downto 0);   -- Registradores de destino (saídas de MEM/WB e EX/MEM do pipeline)
	     forwardA, forwardB		: OUT std_logic_vector(1 downto 0)   -- Saídas indicando os encaminhamentos para as fontes A e B
     );
end Forward;

architecture TypeArchitecture of Forward is
	signal forwardA_interno, forwardB_interno : std_logic_vector(1 downto 0) := "00";   -- Sinais internos que armazenam o encaminhamento

begin
	process(clk)
    begin
        if ((regWriteMEM = '1') and (not(RDMEM = "00000")) and (RDMEM = RSrc1)) then
        	forwardA_interno &lt;= "10";   -- Encaminha o valor do registrador de MEM/WB para a fonte A
        end if;

        if ((regWriteMEM = '1') and (not(RDMEM = "00000")) and (RDMEM = RSrc2)) then
        	forwardB_interno &lt;= "10";   -- Encaminha o valor do registrador de MEM/WB para a fonte B
        end if;

        if ((regWriteWB = '1') and (not(RDWB = "00000")) and (RDWB = RSrc1)) then
        	forwardA_interno &lt;= "01";   -- Encaminha o valor do registrador de WB para a fonte A
        end if;

        if ((regWriteWB = '1') and (not(RDWB = "00000")) and (RDWB = RSrc2)) then
        	forwardB_interno &lt;= "01";   -- Encaminha o valor do registrador de WB para a fonte B
        end if;

    end process;

    forwardA &lt;= forwardA_interno;   -- Atribui o valor do sinal interno forwardA_interno à saída forwardA
    forwardB &lt;= forwardB_interno;   -- Atribui o valor do sinal interno forwardB_interno à saída forwardB
end TypeArchitecture;
</vhdl>
</project>
